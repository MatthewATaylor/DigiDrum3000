`default_nettype none  // prevents system from inferring an undeclared logic (good practice)

module top_level (
    input  wire         clk_100mhz,  //100 MHz onboard clock
    input  wire  [15:0] sw,          //all 16 input slide switches
    input  wire  [ 3:0] btn,         //all four momentary button switches
    output logic [15:0] led,         //16 green output LEDs (located right above switches)
    output logic [ 2:0] rgb0,        //RGB channels of RGB LED0
    output logic [ 2:0] rgb1,        //RGB channels of RGB LED1
    output logic        spkl,        // left line out port
    output logic        spkr         // right line out port
);

  //shut up those rgb LEDs for now (active high):
  assign rgb1 = 0;  //set to 0.
  assign rgb0 = 0;  //set to 0.
  assign led  = sw;

  //have btnd control system reset
  logic sys_rst;
  assign sys_rst = btn[0];

  logic spk_out;
  assign spkl = spk_out;
  assign spkr = spk_out;

  logic        sin_wave;
  logic        square_wave;
  logic        impulse_approx;  // same as square at very high frequency

  logic [31:0] wave_period;
  logic [31:0] wave_frequency;
  logic [31:0] square_count;
  logic        square_state;

  logic        divider_busy;
  logic [31:0] divider_out;
  logic        divider_out_valid;
  divider my_divide (
      .clk(clk_100mhz),
      .rst(sys_rst),
      .dividend(32'd50_000_000),
      .divisor(wave_frequency),
      .data_in_valid(!divider_busy),
      .quotient(divider_out),
      .remainder(),
      .data_out_valid(divider_out_valid),
      .busy(divider_busy)
  );

  always_ff @(posedge clk_100mhz) begin
    wave_frequency <= {27'b0, 1'b1, sw[15:12]} << sw[11:8];
    wave_period <= divider_out_valid ? divider_out : wave_period;
  end

  counter wave_count (
      .clk(clk_100mhz),
      .rst(sys_rst),
      .period(wave_period),
      .count(square_count)
  );

  localparam upscale_factor = 8;

  counter sampled_counter (
      .clk(clk_100mhz),
      .rst(sys_rst),
      .period(100_000_000 / (upscale_factor * 44100)),
      .count(sample_cycle_count)
  );

  logic [15:0] sin_sample;
  logic [15:0] sample_out;
  logic [31:0] sample_cycle_count;

  always_ff @(posedge clk_100mhz) begin
    sample_out <= sw[0] ? sw[15:8] << 8 : sin_sample;
  end

  sin_gen my_sin_gen (
      .clk(clk_100mhz),
      .rst(sys_rst),
      // ideally 2^29 * 2pi * freq / cycles_per_sample
      .delta_angle(wave_frequency << (16 - $clog2(upscale_factor))),
      .get_next_sample(sample_cycle_count == 0),
      .current_sample(sin_sample)
  );

  dlt_sig_dac_2nd_order ds_dac (
      .clk(clk_100mhz),
      .rst(sys_rst),
      .current_sample(sample_out),
      .audio_out(sin_wave)
  );

  always_ff @(posedge clk_100mhz) begin
    square_state <= (square_count == 0) ^ square_state;

    impulse_approx <= square_state && (square_count < 1000);
    square_wave <= square_state;
  end

  always_comb begin
    case (sw[1:0])
      2'b00:   spk_out = square_wave;
      2'b01:   spk_out = impulse_approx;
      default: spk_out = sin_wave;
    endcase
  end

endmodule  // top_level

`default_nettype wire
